module unpacker (
    input [31:0] data,
    output [:0] result
);

endmodule


