module cos (
    input clk, 
    input rst,
    input en,
    input [31:0] x,
    output [31:0] cos 
);




endmodule
