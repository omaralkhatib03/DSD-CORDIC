module fixed2float (
  input [:0] result,
  output [31:0] floatResult
);

 
endmodule
