module engine (
    input logic [31:0] theta,
    output logic [31:0] value
);



    
endmodule