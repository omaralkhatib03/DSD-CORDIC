module iter (
    input [4:0] i,
    input [:0] atan_i, 
    input signed [:0] x_i,
    input signed [:0] y_i, 
    input signed [:0] w_i,
    output signed [:0] x_n,
    output signed [:0] y_n, 
    output [:0] w_n
);
endmodule
