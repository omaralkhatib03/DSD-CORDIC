module controller (
    input logic clk,
    input rst,
    input logic isSpecial, 
    output logic iterator
);


// TODO: Implement controller FSM

endmodule